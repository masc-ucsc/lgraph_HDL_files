module clkGen(clk);
output clk;
reg clk;

initial $clkGen(clk);

endmodule
